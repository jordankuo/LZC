module lzc();
endmodule;